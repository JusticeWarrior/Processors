/*
	Jordan Huffaker
	jhuffak@purdue.edu

	control unit code
*/

// interface
`include "control_unit_if.vh"

module control_unit (
	input wire clk,
	input wire n_rst,
	control_unit_if.cu C
);



endmodule
